`ifndef CONST
`define CONST

`define HV_DIMENSION 2000
`define DISTANCE_WIDTH 14

`define NUM_FOLDS 4
`define AM_NUM_FOLDS 2

`define STOP_FEATURE_WIDTH 4
`define S_FEATURE_WIDTH 4
`define F_FEATURE_WIDTH 5
`define AMP_FEATURE_WIDTH 5
`define FORMANT_FEATURE_WIDTH 11
`define MAX_FEATURE_WIDTH 11
`define TOTAL_FEATURE_WIDTH 40

`define STOP_NUM_FEATURES 11
`define S_NUM_FEATURES 14
`define F_NUM_FEATURES 18
`define AMP_NUM_FEATURES 20
`define FORMANT_NUM_FEATURES 1601

`define NUM_CHANNEL 6
`define HALF_NUM_CHANNEL 3
`define NUM_CHANNEL_WIDTH 3

`define NGRAM_SIZE 20

`define SEED_HV_MSB 5000'b10111110010000100101011000011000010110110101001110001001110111001000000010001111110011111111100101100100101111011101000010110100111111111010101101111101000110111011110100100000101100001001000111010001111011100011001010110010000001110010111110010001001100110101000001001100000001100110000010100011001010101001101001100100110100111101000001000101100110110010000101000010111110000000010100111110010000101011110111101100101110000111101010001110111001101100010000101100110100001000001010010101011011010000010110001100011100011010010101100001000011011101101110110000111110110110111100101001101100011000010001011000010101101110111111110000010011011000101100101011010000001000001111110101010010110001001011010000100001001011000110010110100101010011111100000000010110010011000001000100000111000010100101001100010111101100101100110101100110100101101010001110110100101011010110011001001101000110010000011100111010010111110011001111010110100000001100011110010001101001011100000001110110001111001010001010001000011000011011100011000111001000010010101000110111000001000110100011010111000100100000111100001000011110100100100111110000010000001010111001011010111010110000010111110111111101101010101100111000001101110000000010010000011011010011101011111111100100010010001010011110011101000011101111010101111110101001011100000110110001110010110001111100110100011001000101010101001101111101100000000010011100110100000011011001101000011101111110000101100110011110000011101011101111101011101010111010000111000010011011110010100011000011110011101110111111011010000011101000001011011011010111101000000000101110000100110001111110111101100010101100100110110100001010010100011100111111111011001111101110101111111101010010000100111000000100001011101011110110000101100011001000010011011000000101100001110010100001110001110101000101011010010001010011110000100101101010101010001010100001001100101100000100100001001000110100011010011000100100111001101110010100110011110001100101001001011100011000111100001000100111101101000011001100101000100001100010100011001110101001101100001101100011000010111001111011110100000011100100010100000111011001011111101111101000001011001101110001111010001110110101000000000101111101100010101000101111100110101001111001010111101100000011000101101010101101011010101011110110010111101011000101011110100001101100100110001110101011001000101000111111000110000011011101100001100000100000101001011111001000101011100000010000001110100000101010111011111110111011111111101001010001000001010101000111111111100001111101110110100001100101011110010111111000100001100110111111010100010110010111001011010100100000110000101110001111010111011010101000101101110011010011100100100001100111010001101001010010110010000100111001011110100110100000011111001011000111111010000100000000011110100101101111101100001111101110000101001110001111010011100100000011000010111001100010101000111101010011001110101100101001001110100000101011101100010111011101101110101011111001010010101010000010101011101101000011010111010000101010000010101111011000111111100100101110101101000100111100110100000001011110000011111010111110110101111010011010010000100000101010101110001011000010110000000100010101110101000110111001000101100011000111010101010000000111100110000101011101010001001110011001000011001111111000011111110001111011111101111100100001000111011101101100011001101111001011010101010001100010000011000111110111011111010010100101000001010110101110000011101100100011110000000100100111011100010000111011100111111100001101101010011000011010001001101100000001111101101111110011001101101000100011010110001111100011001010110001000000101111010001110100011101100001111101011111110001101000101001001010100010101010111010000000101101000010100010111110110001010010101100100100111100101010010111011101000111110011110101110011011110010111111111011001010011111111110001000000001001001010000001101110101000001110100111001001001100110011110000110111110011010111100101110100101000110111110111001100111001010000010001001100011111111001110101010110011111001101001111001100100010100010100100011001100111001110010011011101110011110000010101110001101010001011010110111111010011011100110110101001001001101111110101001000100001100001000010110111100001110011100011101011010110100001111011001011010010000101011010101101001111100010101111000110010101011110110100100011110111000000110000011110110001001011100011001111111011000001001110110001011101001000001000000001101010010000110010000101001110011110101001110100100100111111000101100011100001110000001000000101011111011001101110100000100110101100110100011001000000110010100110100111000010010100010010000010010010010101011000110100111101001011111110001010111000011010001010101110101000010000011011110010101011101011111110100110000011110001110001101011010011000001011111101001111010101100100010001000100100111110100111000110010111001001100010110111111001010011001101100100100011010101100000000101011110000010010101100100111111010111000001001000010010011010101110100000010011010111100011100010001111100110010111011110111001
`define SEED_HV_LSB 5000'b00110111101100010000000111101001111111010100000101110111100010011111011011001010101010011111000001000110010001101100100111001010101011001000100101100111001000001110111101110100010111100100011101110011011010110101011101101101001110010111111100110101010111111010000110111011100011101000100001011101100010000101011001010010000100010100111110001001110001000111001010100010110001001000010010101000000100111111011110101101101101001011100100010111101111100101010111000111010101100001000110111100010001011000001100110011111110111000111111100001000010110000110110110111010101011111110110011000101100010010110100101011100100100000111110010010100011110100001011000011101110011001001011100101101101000111101110010101111011101101110111111101100000100001011111010100000000101001111111000001110101010010011001000010111011110000111010110100111111011010100101101110010011100111101011001111000100010111101011101001001010000101111111000011101101101101101010010010001101011011101010110001111110001100101011010010011111101110010101101101100110001101011110101000100111010001011100011101100111111011110000111110111100110110001001101010100111011001010111110111100011100000100101100001001101101111010111010001011010011100100011010111010100101010001000110100101011011111110111011000111110001101111101001011011111101101110010111110010010111001101001101000010101000011110110001011110000010001101110010111001100101110110100111000110101011000100001000101111100101100010000010011101010111001000101100001100110100000011110110011101011101010101010111100001100001101001110110100111000001101111101001010010000011000010000110101000010100100010001111001101111001100100001111111110110000010111011000110111000001100011101011010010001011011011010000011010111001100001110011000010010100111101011101111111100111110011100000011111010001000111001000101101110110110100011101111101111100100010110010101001111101111001001100001111010011110000111110101100011110011000000001101011011010001111000110100001110011011100100010100000011001011010001111011010100001101011101110000011100000110011010010101111111111010000000110111110101110000011010010101101110111001000011110010111010000010101000111011111110000111101101000001110001010101100110000001010110011111100100100101101101011011001011000101110001111001001010000100100011111000110011100001100101011101010001000101011110101111011101110010100101010010111011001011010000100011100111110000000101110101001010100101100111100000001100101100001011010101010011100100100101101000110011011001001001110000010001100100011010111110100100111010101111110001000101100110100010100110001111101100010000001000100001110111001100111001000000101110111111110010010000111100110110101111010011111101101001010011101101100011100011010100000001111101111111101001000111101111010000100011100100111110000011011111100101000000111001011100111010011011000000110101111000110001110111011010111011010101110111101010101010111111010000101011100000001111101001101011111011110001011111000111010011111111010001001110011101100111010001101101000100110111100010110100011000101011101001100100001110110011000000010010110000011011101100000111010111010011000110001101001000100000110001000110000001111011010100111010100111101101010101011111111100110110010010100000011001000101110010010010000011000111001000111111011011100010010100010101000100000111110011101110101000100110000011110111110000011001000000011101111010111010101001011001110110101001000000011001101111001111100110001101001101101001000011110001100101100001100000000101111110010111110000001110011100001111000100111011101111000000011011111000010111100010110001110011110110001000110000101010100110100101001011001101010110100001001100001111010001110001100000110100111010101100011000001011000001010110000111011010000100011111101010000010001000001100110101001010010011010000101001100100000101011101110110000100000110101010101110000101011101010011000001011010011101101101001110100110001111010111000100110011000111000111100001101110001110001111100001101000110000000011111010001101111111110010110011010011110001010011011001100110001101010111111001010111000010111011010000101111000111010111000000011110001000110110001011110101110000110100110110101101011000101000011100101010001101100100001011100110000011100010100000111000100011100110001000011010010100001011111100001010010001110111001000111110000001110100001110010101011001000000001001010000010011100110010101000011110001010101101011111100100001001010001111101111001111010111110001000001011011110010111111001000111101001110011001101110110100101111100001111111111010111100100010100110111101100011001001111111011000010000101010101100001101000011110111001010111110110100110011001101111100001001000101011000100000101100111011101011000001111110101100101100011101000101101100001100100110011101101111101110001101010001000010110001101111101011111101010111100100000011000111111000100011100000000101101001101011000101110000111111000110111010100010111101010111111011011001110000111100000010110001010001100001000000001000111101100110011000111010101111001100100110


`define ceilLog2(x) ( \
(x) > 2**30 ? 31 : \
(x) > 2**29 ? 30 : \
(x) > 2**28 ? 29 : \
(x) > 2**27 ? 28 : \
(x) > 2**26 ? 27 : \
(x) > 2**25 ? 26 : \
(x) > 2**24 ? 25 : \
(x) > 2**23 ? 24 : \
(x) > 2**22 ? 23 : \
(x) > 2**21 ? 22 : \
(x) > 2**20 ? 21 : \
(x) > 2**19 ? 20 : \
(x) > 2**18 ? 19 : \
(x) > 2**17 ? 18 : \
(x) > 2**16 ? 17 : \
(x) > 2**15 ? 16 : \
(x) > 2**14 ? 15 : \
(x) > 2**13 ? 14 : \
(x) > 2**12 ? 13 : \
(x) > 2**11 ? 12 : \
(x) > 2**10 ? 11 : \
(x) > 2**9 ? 10 : \
(x) > 2**8 ? 9 : \
(x) > 2**7 ? 8 : \
(x) > 2**6 ? 7 : \
(x) > 2**5 ? 6 : \
(x) > 2**4 ? 5 : \
(x) > 2**3 ? 4 : \
(x) > 2**2 ? 3 : \
(x) > 2**1 ? 2 : \
(x) > 2**0 ? 1 : 0)

`endif