`include "const.vh"

module associative_memory #(
    parameter AM_NUM_FOLDS, 
	parameter AM_NUM_FOLDS_WIDTH, 
	parameter AM_FOLD_WIDTH    
) (
    input                       clk,
    input                       rst,

    input                       hvin_valid,
    output                      hvin_ready,
    input  [`HV_DIMENSION-1:0]  hvin,

    output                      dout_valid,
    input                       dout_ready,
    output reg [3:0]            keyword
);

    reg  [AM_FOLD_WIDTH-1:0]        similarity_hv;
    reg  [`DISTANCE_WIDTH-1:0]      distance_ON;
    reg  [`DISTANCE_WIDTH-1:0]      distance_OFF;
    reg  [`DISTANCE_WIDTH-1:0]      distance_GO;
    reg  [`DISTANCE_WIDTH-1:0]      distance_STOP;
    reg  [`DISTANCE_WIDTH-1:0]      distance_LEFT;
    reg  [`DISTANCE_WIDTH-1:0]      distance_RIGHT;
    reg  [`DISTANCE_WIDTH-1:0]      distance_YES;
    reg  [`DISTANCE_WIDTH-1:0]      distance_NO;
    reg  [`DISTANCE_WIDTH-1:0]      distance_UP;    
    reg  [`DISTANCE_WIDTH-1:0]      distance_DOWN;    
    wire [`DISTANCE_WIDTH-1:0]      distance;
    reg  [`DISTANCE_WIDTH-1:0]      curr_min;
    
    wire                            hvin_fire;
    wire                            dout_fire;

    reg  [AM_NUM_FOLDS_WIDTH-1:0]   fold_counter;
    reg  [3:0]                      prototype_counter;

localparam PROTOTYPE_ON = 10000'b0111000011111000010001010011111111100001000001111111000100111100101100001111000011100011010001010100110111111010111000110101110011011110010000011100001000001100010111100010100001110110000110010111010111110101101111101111101100101000011101111110001110010001110001110000111110001100010011101000100000000010001100001100110101000011100001001100011101111111101101000010011101011110011011100000100100000110101100111001001101001000101000011000000011011100110001101101001100101100011101011011100010111111110010111111001000000000001111101010111011001110010010111110000010010010101000001101110011000000100011001000101101010111100011111111100010100101111010001111010111110111100011100011010101100001000011001001000100011010101011110000111100101110011101000001011100101111110011111110000000011010011101110110000110000011100010100000111101110110000110100100110011100100110011001110000001000010000111100111001001100011111000010111100111001100101000100011011100000111000111110001110110001001010100101000110011000000101001100001110011111000110011100001101111111011000000101000110010110000111101110011000000000111111000011111110101100100111000011101000110111000101010001110010000101110010110111111101101000000110111100000000110100100001111000111010011000111110010111100001111000001100000010001110111000010001111111110010100100000000111011110001000011101100001100111111011011111101100101001011010100101001010010011011001111100101010000001011111000111010010000111111001100100111101001000100001110111001011001111011010010010111110011110011000110011001100010110010010110111111000110001111101100110101011101011100100000110000011010110001000101100010000011111011101010100100101000111011000100110111111111110111111110111011110001110010101011111111110100110001111000000111111011111110100000110101001111111100101110001010101101110011100000110011101110000100110001101101100110010100001000100011110001101001111100111111001100011101111111110010100000111111111100001110000001100111111011110110000000110101101011100011110011000101010010000011100101101101010100110110100110010111101011010101101101111110100010001010110101101000000001010100000000000010011111001111011011001100010100000101001110000011011110111100001000110101000011111010000000110110000001001111011100110001101011100001110100111001000011111010110110110110100010011001110010011101000101010110000000101010010001110001111111001101100000101000000011110000000000111100011110011110000111111010001110011001001011111001011010110000100100001000000101000100000010011111101100111101111010000111101111000011110011010100010000011111001000101011101011101100011101110101100110000011011101010001010000001100001001111101011110110010001010111101000110010010000111011111100011011100011000111101100111001010111010001111100111110110011100000001001111100000111010100100111111111110001000000011110111101001011110000010110000111111000101010011001101111100000000001000101010001000011011011101011101100100111101010011101001010110011001111010011110101100110110101001100010111100111001101000011001111100000100111101111111111011001100001010011110000000001101100001010010100100010011100111111100101010001110001001101011000000111001110001000000000100011100111001110010011101000000111010110001101100110000000101101110110010001000001101010110011101101000100110001001000110101001101000111110001000101010110011011100010011001000111111000100111100001110000010101011000100011011111110010100011001110011000110011110111010100100001101101100100010101110001011001010000011110001111111000001101010010000000100011010110101111010011011101011110101000100010100100001001111011110000001111011100101001010100001011001000011100000011011010011110000011110110001110000101101100100001111110011011110000101001000000000000001000111111110101000000010000001010100100011001111010000001000011011111011000000111100111110001011110110001000100100000111110000000100000110111101111111000110010100100000111110011111010001011110111010101010000101011111010001000001100000011011011000101010100110110010110100000110101011001011100111101110001010001100010011001010000001011011101111101111101010001101101011110110010000101000010100111010101000011000001010001011110000010101111110110100000011000111010001000000111101000110001001000110000111100010011110110110001111101001011001010011100111011000011010100101000101101100100010010110100000101000001101010110010001100011111011111100111011010010000100010110001011000000000111111000010100000000001110000111101110110010001110001100010111001110010111010011011000010001101100100000000111111000001010001011011001010111101110111011010100000001110011010100100100100010100010110000010000011010110011100001101110001000111111111101100101111001000011001111100101011000011011101011000100111100110111011010001010000100111011101111011111100011110000001000001110000100100110011010000100100000000000011000101000000011110001001110101010011111101100100011000011010000010110000001000010011000111111011110000001110010000100001100000010011111101110010000001100010110000100011110010000101111011001000101110010010101010110111111011111000010011110111111110001100111001111101000010001101101111010010100010100100001001101000011111000100010110001100100101110000000011110000011001110111000001111100110001110010111001111101111101010010010111100001011000111101110110000101000100000011101100010101010111011100001110100111111001011010110110101010001001010001111111110001101101100110000010001011100101011011110011111100000000110101100011110011110011011000110011000010000011101110001000000000110110000000011111110101100110110000001111000101110111110000101110010111011111010010000100000100011111000001100100111110000110010011111100010010001100110111000000111111111110011111100010000111111100010110100111001101011111010001101011011100001000000011001111000110011101011110011100000001001000011000110111001001110000101000110110011101001000110010110011001111100101000100001110000110100000101100010011010101000011111101100111100101011111100110110110011111100001010110110100010011000011110110110110011110001110101100101001001011110110000100000000000000111100111101011011110001001100001101011100001100001101000001110000110111011111100011101011001001000110000110011110110001100000000000010001111111000110011000011110100011001110010011101011001011011010001101100010000001011001000100111000001111101001111000000110111000101110001111111001110101111111011010010000011010111100111011111001101110011100111100110011010000111110110010001100011111001101010011111000011111111011001111011100010000001000110101011000000101000111011100100011011001101000110110100011000101010010011010110001101101001011010111100110001001111111000100001111000100101100011011101001111101011000010111111110100101011001111110000100000101101100111011100011111111110011000000110000111100000100001101001010010110110100110100111100111111010011000001010011001111101000111100000000111101100000111010101100110100110000001100001101001101001111111000100111100100001101001111001001000000111001111110111100011001000111010000000101110010100001001101101110101111000100100011000110010111001000010111111011100101110110100011011100011100000111001110000000101000001101110000100101100100100001110010001000011010000110001000101001010011100001101101010001110001100010011000001111010110001101001111000011111001110111111001001110100100000110101111111101111000100011110011011100011001000100011100111010000110000011111100010100001101101110110101110000101001110111011100110110100111110000000010111111100001100101000011111001011110010101111011100000011000100101100110110110100110110011001110000100011100011101000000001011010111111110111000010000110000011000010110011111000111011110000110100101100111000010110110000001001110101010111000010011011101011010111100110011110110011000110000011101101110000000011100000101011011001101001000111110000000010000100010111001000001001111101101101011010101001011100001000101100000111011110100111100101110000101001001110101101110001111010001000010001111000101100101101110000000011001100000111001010111011011011100100100001110110111011001100101100111000000010010110101001000110011000100110011111011100100110111111100001011110000001001001100001011101100011110000000001110101001010110011000000111010110011001111100001100001111011011100010001110000110010011100001100100001101111010100001100110111001001110111110000011101111111001101010111000010001111110111001011001111101111000010011100000010110001011111110010010111101000011011100001110111100011010011110010111011101101100111010001001110011110100000100100110000111011000000000010000110101101000111100110100111111110000000011111000100101010110000001101010111011100010001110111111111011010010110111111010100100101000001111010100001001110111011010010011010000000001001001110101010100110001100110111111100011000000110110110001011011111100100111011010101011001111011101111010001010100100110110101010001010010110100000011000000111110100000001011100111110010101100101110001000110010000000110101111111110001000111111010001111100100001110011000001011000000011000100110111111000000101100110000100011000100110111111101000100000001010111011110011101111100111000111011011000110000001000010011110100111000010011100100100000111000111100001111101000000010111100001000010000010011000001001010110011111000000100111001111111011011101100010000110111000000100111000010000110101101111101110001111000000100100111011010001000011111011011111111100010001011101101100000111011001010010000111011001101111100000010110011101110000000110101000111101010101010001100101001001111011000000000001001000001000010001000001101110010001010001011001111000101001001010011011110100100101001111111111011100110001000000110100110000101100110011001110011111001100110111001000101011110111110111100100011110111000000000001111000111000000111100001110101111010101101011011000110110011000111100110001101000000111011100011100100010000000110000010001110010010110000010001000110011001110010000011111011110010010011000001110100000010000000111100111101111000100000001100000010000010011101001111001101011110011000001011110000010001000000001111100010001111010100110100001101110;
localparam PROTOTYPE_OFF = 10000'b0110000011111000010010110010111101100011000001111111000100110100101111000100001011101011000001001100110001111010111000110111110011011110010000011100000110001111000111100010100010110110000100000110010101100101101111101111101100011111001101111110001110010011110001110000111100001100010011111000000000100001101100001100110001111011100000101100011111111110001110010010000000111110011011100000100100110110011100111001001101000000100000011000000011000100110001101101001100101000011101111011100010011001110001111111001000101000011111101000111011001110000010111110000011010010101000001101110011001000000000001100101101100101100011110111100010100101111010001110110001100111100011100001010101100001000011001001000100010111001011110010111101101110001100100001111100101111110011111110000000011011011101110110000100000111100011001000111111001101000111100100110010100100110010001110000001010011001111100111001001100011100000010111100111001100101000100010111100010111111100101111110110001001110010101000110010001100101001000001110011111100110011100001101110011011000000101100110010110000111101110011000011110101111000011111100100010000111000011101000110111101101010001101010000011110100110111011110001010100110111100000000110100100001000111001000011000101110010001100001110000001100001010001110001000010001111111110010110000000000111011110001000011101110101100011111011011111101100101001011001100101010010100011011001111100101010000001011111000111110010000111111001100100111101001000100001110011001011001111000010010010111110011110011011111011011110011110010010011111111100111001110001100110101010000011100100000110000011010111111000101100001000011111010011000100100101000111010100100100011111111110001110010110111100000110000101011111111011100110001111000000111111111111110100000110001001111111100110010001010101101110011100000110010111110000000110001100101011111010101101011000011100001101001111101011111001100011101111111110010100001111111111100111111000000110001111011110101110010101001101011100011110011100110010010000111100101001101010101110111100110010001110011010101101111110110100010001010110101101000110001010100000000000010011111001110001011001000010100000101101110000011011110101100001001100100000011111010011000110110000001001111011100110001100001000111110100111101000011111010110110110110101010011111110000111101000101010110011000111010010010010110101111000100000000110000001100010010111100111100011110011110000111101000001110111001001011011001011010101100100100001000000101000100001010000001101111011101110010000110011111001011110111010100010000011111001000100011010011101100011101110101100110000011011101010000110000001011001001111101011110110010001011111101000010010010100111011011100111110100111000111010110110010010011010001111100111110110011100010001001111100100111110000100110101110010111000000011110111101001011000000010011000111111000101010111001101111100000111010000001010001010110011011101010000010000111101101011100001100100111111111010011110101100111110111001100010101101111111101000011101111000000100111001011110111011001100010010010111100000001101100001010010100100010011100111111010101010001110001001101011000001111000010111001000000100010110100001110100111111010000111010110000000110110000010101100110010001111000001101010010011101111000100110010001000010101001001000111110001000101110100011011100010011001000111111001010111100001110000011101001101100011011111010010100010001110011010001011110000010100100001101101100100010001110001011001010000011110001111111000001101010010000000100011010110101001010010000100100010100000100010100100001010001011110000001111011100111001010100010011101010110100000011011010011110000011110011001110000101101100111101111100101010000001101011000000000000001000111111110101000000010000001010000111011001011010000001000011011111011000000100110111111001000000101100000100000100111110000000100000110111101111101000110010100100000111110011111010001011010111010101010000101011111000001001001100000011011011000101110100000100010110110000111100110101011100111101110001000001100010011001011000000011011101111101111101010001001101010000110010110100100000000111010100001011001101010001011111000000101111110110101100011000111010001000000111101000010001101000110001111100010011110101110000000001001011001110011100111011000111010100100000101100111000010010110100000111001001101010110010011101111111010011111111010101100111100001110001011000000000100111111110100000000001110000111101110111010000111001100010101001110000111011011011000010001101100100000000111111000001010001011011001010111101110111001010100000000110011010100110100100010101010110000010000010010110011100001101010001000001111111101100000111010000010011101100110010110011011101011000011010011110111011010001010000110111011011111011110100011110010001000001110000100100110001010000100100110000001001000101000000011110011111110101010011111100011101011000011010000110100000001001100011000111111011110100001111010000100001100000010011111101110010000011100010110000000000000010100101111010101000001110010010101010110111111011111000010010010111111000111100111011011101000010101101100111010011100011000100001001101001101011000100010110001100100101110000000011110000011010110111010001100100010001110010110001111101111010010010000111100001010011111101110001100101000000000011101100001010110111011001101110111110111000100011101110101010011001010001111111110001101101100110000010001011100100111011110010000000000100110100100011110011110011011000110011000000000011011111111000000000100110000001111111110101101001100000000111000101010111110011001100100110011111011000000101110100011111010001100001111110000110101011000000010010001000110011000000111111111110011111100010000111111000110110100111001101011111110001101011011001111000000011111111000001011101000010111100010000001000011000111111001001000000101000111000010101110110110010110011001111100101000110001110001111100000101100010011000101100011111101100111000101011111100110110110011111100001010110100100011000000011110110110100011110001110101100101001010011110100000100000100000000111110111011101011111001101100001101011100001100001101010001100001111111011000000100001011000101001010000010011110000001100010000000010001111111000110011000011110101011001110010011101011001011011010111101100010000110011001010100111000001100001001111110000110111000101110001101111001110101110101011010010000011010001101111001111000011110011100111100110011001100111110110011001100111111001101010011101000011111111011001101011100010000001000110101011000000101000111011100100011000001001000110110100111000101010010011010110001101101001011010111100111001001111111000100001001100100000010001111101110111101011000010111111110100101111000011110000000000100001100011011100111111111110011000000110000111100000100001010001011110110100100110100111101001111010011000001010011001101101000111100000000111101100000011011001100101100110000001100011101001101001111111011100111100100111010100000000001000001111110000010111100011001011110010000011001110010010001001101101110101111000011100011000110010111001100010110011011100101110110100000100100001110100111001110000000101000001101110000101110011100000101011111001000011010001110001000101001010011100001101101010001110001100110011000001111010110001101101111000011111001110111111001011110100100000110101111111101111001111110110000111101010001000100011100110000000110000011000100100011001101101110110101010010101001110111111110110110100111110010000010111101100001100010000011111001001000010101011011100000011000111001100110000110100110110011000110000100011100011101000000000001010101011111011010010111110000111000010110010111000111011110000110100101100111000010010100100101001110001010100010111011011101011010111100100011110110011000110000011101101110000110011101000101011011011101001000111110001000010000100001111001001011000011101101100000100101001100010001100101100000111011110100111100101110000101001000011011100000001110110001000010001110000101100101111101110000011101100000111001010111011011011010110110001110110111011001100101100111000000010000010101001000111011000100110011111000100100110111111100001011111100001100101100001010101100011110100000001110000000000110011001000111010110011011111100000001111111011101110000001100000110111000100001100100001001111100100001100110101001000110111111100011101111111010101010111000011001111010111001011001111101111000010011100000010010001011111110010010111101000011010110001100110100011010011110010111011101101111001010001001110111110100000101000110000111011000000000010000110101101000011100110000111111110000000011111011100101010100000000101010111010101100001110011111101011010000010111111010100100101000000111010011000110000110111010010011010000000001100000010101110100011001101001011101100001110000110011110011111010111100100111011010100011001111011101111010001010100100110110101010001010010110100000011000000111110100000001011101111110010111100001001001001111000100000110001111111010001100111111010001101100000001110001000001011000000000000100110111111000001001100110000100011000100110111101101000100000001010111011110011101111100111000111011011000110000001000110111110100111000010011100100100000111110111100001001101000000010111100001000111000010011000001001010110011111000000100111000011111011011101100000000110011000000100111000000000110101101111101011101111000000100100111011010001000011111011100001111101010001111101101100000111011001010010000111011111100110010000010110011101110000000100101000111101010101110001100001001100101010000000000001001000001000010001000001101111100001010001011001100000101001001010001011110100100101001111111111011100110001000000000100111000110010110011100111011111001100110111100000111001110111110111100100011110111010000010001111000111000000110000001110111111010001001010010000110110011000101100110001101000001011011100011110100010101101011000010001110010110110000010001000110011001111010000011111010000011010011000001110111000010000100111100111100101101100000001100000010000010001101001111001101011011011000011011101000000001000000001111110010011111000101000111000101111;
localparam PROTOTYPE_STOP = 10000'b0110000011111000011110111100111111100001000001111111000100110100101111110100000011001011010000111100110011111010111010110101110011011110010000011100000110001111000111100010100000111000000110010111010111111101010001101001101000011010110101111110001110010001110001110000111000001100010011111000000000000001101100000100110101100011100000101100011100000000001000000010011101011110011011100000100100110110011100110001001101000000100000011000111010011010110001101100101100100100010101111011100010011000011010110111001000100000100111110110011011001111010010111110000011010010101000001101110011001000100100111000101111011011101011111111101001100101100110001101010001100111100011100001010001100001000011001001000100111101011011110001011100101010101011000001011100101111110011111110000011011111011101110110000100000111101001001010111111011101111110110111110100100000100011001110000001110011001011100111001111101011000010001011100111001100101000100011010101000111000111110111110110001001000010011100111101100100101001101110000011111110110011100001101100111011000000101000110010110000111101110011000000000111111000011111110100010000111000011101000110111000101010001100010000011111011110111011110001011100000001100000000010100100001111111110010111011001110010111100001111000001100001000001110001000011001111111000010100010000000111011110001000011111110001011011111011111111101100101001111010000111010010010000011001111100101110010001011111001110110010000111111001100100111101001000100001100110001011001110000010100010111110011110011001111011011110010110010010111010111000101001111101100111011100010111100100000110000011010110001000101100011000011111011101000100100101001111011000100100011111111110001110010111011110001110010111011111110101100011001111000000111110010111110100000000001001111110100101110001010101101110011100000110000110010011100110001100101100111010101101011011011110001101001111101011111001110011101111111110010100101111111111100101000000000010000111011110110000000110101101011100110001100100110010000000111100110101101010100110111100010010111101011010101011101110110100010001010110101101000111001001000000000000010011101011110001011001001010100000101001110000011011111000000011011000101000000111010010000110110000000000111011100010001100000001001010111011010001011101110110110110110111010011111110010011101000101010110000001110110110001000001101011001100000001111000000011110000110100111100011110011110000111110101001110011100000011011001011010100100100100001000000101000100000010110001101100011100110111000000011011111011111101010100010000011111001000101010001011101100011101110101100110000011111101010000110000001100011001111101011110110010001011111101000010010010000111011111100000001111011111000011010110001110111010001111100111110110111000000000001111111100111010111000110100110010111000000011110111101001011000100010011000111011000101010001010011111100000000000000101000001010111011011101011000000010111100101101101101100110101111011110011110101100111110111001000010111110110001111000011101111000000100111101111110111011001100011010001101100000001101100000110010100100010011100111111100100010111100001000001010000001100101110111000000000100011100100001110011011101001110111110110111000111110000010101100110110001111000001101010010100010011000000110110001000010101001011010011110001000101110100011011100010011001000111111001000111100001101000010101000100110011011111110010100010001100010010110111110110001100100001101101100100010010001001011001010000011110101111111000001101010010000000000011011000100111010011000010100010101000100010100100001110001011110000011011011100111001010100010011101010110100000011011010011110000011111000001110000011001100111101111111100001000101101011000000011000011000111110010101000100010000001000000101000101011010000010110011111111011010000100000111110011001000101000011000000000111110101010100000110111101111101000110010100100000111110011111000001011001111010001011000000101111010001000001100000000000111000101000100000110010110100000111100110100011100111101110001010001100010011001010000000011011101111101111101010001001101010001010010110100100011100111010101000111001101010001011110100000101111110110100000011000111010001000000111001011010001101000110001111100010010111101110000111101001011001110011100111011000111010100101000101101111000010010110100000110001011000110110010011101111101011111111111011000100000001010101001001010000000110111010010100001011101110100111101101110010000111001100000100001110000111011011011011010001101100100000000000111000000000001101000101010111101110101011010000000000110011000100101100100010101010110000010000011011110011100001101100001000111111111101100101111011000010001111100101000110011011101011000011010100000111011010001010000101110100011001011111100011110011101000001110000011111110001010000100100111000000011000111000100001110001111110101010011111101100100111000011010000010101000000001100011000111111011101100001110001000111001100000010011111101110010000111100010111011000100000010000101111101000100001110010010111010100111111011111000110010110111111000011111111011011101000010001101101111010010100010100100001001101101100011000100010101100000110101110000000001110000011111110111000001100101110001110010111001011111011010000010000111100001001000101101110001111101110100000011100000010101110111100101000110100111111001011010111110101010011001010001111111110001101101100110000010001011100101011111110010000000000000110100100011110011110011111000110011000000000011111111111000000000100001000000111111110101101000101000000111000101100111000001001110010110011111101000000100100100011111010001100001111100000110010000100000010010001000110001000000111111111111011111100010111111111100011010100111001101011111101111101011010100000100000011110111000001011101000010100010011000101000011000101111001001110000101000010100110100110110011010110011001111110101000100001110001111100000001100111111001001100011111101100111000101000001100110110110011111100000011111011010011000000100000110110110011111101110101100100111001011110110000100000000000000111100111111001011110001100100010001011100101100001101011001100000111110011101100100001011001010011111100010011110000001011110000001010001111111000110011000011110101011001110010011000001001011011010001101100011110111011001110100111000101100001001111001000110111000101110001001111001111101111101000110010000000010001101111011111111101110011100111100110010001100101110110011101100111111001101010011111000011111101011001001011100010000001001110001011000000101000111011100100001011001101000110110100011000110110011011101001111101101001010110111000111001001111111000111101111000100100000001111101110111101011000010111111110100101011001111110011000000100000101101011100011111111110011000000110000000010000100001101101011110110110100110100111101001101010011000001001011001101101000111100000000111101101000010010101100101100110000001100011101001101001001111011100111100100000010001111000001000000111110111000101100011001010111001100111101110010010001001101101110101111000100100001110110010111001000100100000011100101110110100001001100001110000111000110000000101000000101110011111111011100000110101010001000011010000110001000101001010011100001101101010001111101101010000001101111010110001101001111000011111001110111111001110000100100010110011111111101111000111110110010111101010111000000011100111000100110000011001100010011000101101110110101010000101001110111101101110110100111110010101110111111100101100001000011111111100000010111010111100000011000111001100110110110100110010001010110000100011100011101100000001100110101010000110110010001111000111000001010011111000111011110000110100111100111000010010110000101001101011010111000010011011101010110001010001111110110011001110000011101101110000000011101000101011011001001001000111001111000010000100010111001000001001111101100000111100111001111100001000101100000111011110100111100101111001010101011111011000000001111010001000010001110000101100101111101010000011001100000111001010110011011011010110100001010110111011001100101100111000000010010010101001000010001000000100011111000100100110111111100001011110000001101001100001011101100011010100000001110101001010110011000000111110011011010111110000001111111011101110001001110000110110011100001100110001001111100100101100101001000000000111110101110011111011100101010111000010010100110111001011001111101111000010001100011100010101011111110001010111101000001011101010000111100011010001110010111011100001111001110001001110111110100111111011001100111011000000000010000110101101000111100110000111111110000000011111011100101000100000001101011000101100000001010111111101011010000010111111001100100111010000110000101001101110000110010010011010000000001001101100111010100011001100010101101100001110000110110110011011111111101100100101000011011001111011101111100001110100100110110101010001010010110100001100100000111000100000001011100110010010101100101110110001111010100000010001111111110001000111111010001101100010001010001000001011011001010000100110111111000001101100111100100000000011110111101110111100000001010111011110011101111100111000101111000000110000001000110111110100111000010011110100111100111000111110001111101000000010111111111000011110010011111001000010000011111000000100101001111111011011101100000000110011001000101111000000000001101101111101110010111001000100100111011010001000010111111101101111101010001110101101100000111011000100010000111010001100110010000010110011101110000000100101000111101010101001000011111001000101011000100000001001000001000010011100010101001110001100001011001111000101001001010011001110100010101001100111111011011000000000000001000011100110011110011100001011111101100110111001000111101110111110111100100011110111010000010011111000111001000110100001110001111010001101011101000110110011000101110000001101000001011001111101110110010100000011110011111110010010110000010001010001011001111001100011111001110011010011010001110111000010000011110100110101110101010000001100000010000001111101001111001101011110011000001000111010100001000000001111111011011111010101110111010101110;
localparam PROTOTYPE_GO = 10000'b0111000110001000010001010000111111100001001001111111000110111100101000010100001011101011010000111100000001111010111010110010001111011110110000010100000000001111000111100010100010110110000110010001110011111101111111101100010000101000111101001110001110010001110001110000111000001010010011101000100000000001101100001100111101000011000000101100011100000111101110000010111101001110011011100000100100110110101100111001001101000000010000010000000010011010110001101101001100100011001101011011100010011111110010111111001000000000000111010110011011001110100010111110001101110010101000001101110011000111111100111000010010011010011010011111100010100101111010001111010111110111100011100011010101100001100011001001000100111110101011010010111100100110011100100001101100101111110011111110011111011111011101110110000110000111101011000000111101110101111111110111010011100101110011000110000001100011101011100111001111100011100000010111100111001100010011100011000001000111111011101111110110001000000010011101101101100000101001001111000011111110110011100001101101111011000000101000110010110000111101110011000011110111111000011111110101100100111000011101000110111000101010001110110000011111101110111011110001010010110111100100000110110000010000111001011111000111110010111100001111000001100010011101110001000011001111111110010100011000000111011110001001011111110001011011111011011111101100101001011010111011110010010000011001111100101010000001011111000111110011000111111001100100111101001000100001101100000101101110000010100010111110011001100010110011000100010110010010011001111000101001111101100111011110101011100100000100000011010110001000101100011000011110011101000100100101000111011000100001011111111110001110010111011110001110110111011111110111000101001111000000111110011111110100000111101000111110100101110001010001110110011100000110000011110011111001110101101100110100100001000100011100001101001111100111111001100011101111111110010000100111111111100000010000000010000111011110110010000110101101011100110001100100101010000001100100110101101010100110000100110010001101011010101101011110110100010001010110101101000111001010000000000000010011111011100011011001001010100110101101110000011011110110000011011100101000000110010000000110000000001001111011100110001100000011011110111011010111011101110110110110110100010011001010010011101000101010110011100110110010011110000101111001100000001101001000011110000000100111100011110011110000111110101001110111100001011111001011010110000100100001000000101000100000010001111101100111100110010000000011000111011110010010100010000011111001000100011010011101100011110000101100110000011011101010001010000001100001001111101011100110010001011111101000010010010000101011111100000001110011111111101110110010110111010001110000111110110011101100000001111100000111010000100111111110010111000000011110111101001011000000010111000111111000101010000001101111100010011010000001010001000100111011101001001100010111100101011100001101100011111000110011110101111110110101001100010111100110000001000011101111000000100000001011110100001001100001110010110000000001101100001110010000010010011100111111011100110111100001110001010000001111101110111000000001011110110100001101011000101001111011010110110010010110000101001100110110001111000001101010010011101101000000110100001000010101001101111011110001000101010110011011100010011001000111111001000111100001110000111101000100100011011111010010100011001100100110100011110011010100100001101101100100011010001001011110010000011110001111111000001101010100000000100011010100100001010011000010100010101000000010111100001110001011110000001101011100101001010100110011001000110100000011010110111110000011110001001110000111001100111001111100000010110101101011000000000000011000111111110101000000010000101010000100011001111010000001000011111111011000000111000111111001000110011110000100000100111110000000110000110111101111111000110001010100000111110011111010001011010111010101011000000101111010001001001100000001000001000101001100000000010110110000001001111010111100111101110001010001100010011001011000001011011101110101111101110001001000010101110010110101000010011000110111100011000001010000001111110111101111110110111111100010111010001000000111101000110001000000010010111100010010111101110001111101001011001110011100100111000111010100100000110001111000010010110100000111000001101010110010011101111001011110000111011010110111100000110101011000000000111111000010100000011001110100111101110111101001111011100010111001110000111011011011011010000100100100000000111111000000010001101000101010111101110101010001000000000110011010100100100100000100000110100011001011011110011100001101110001000111111111101100101110110011110001111100010011000011011101011100100111100010111011010001011110110111010011111011111100011110000001000001110000000111110001010000100101001101001011000101000000010010001001110101010000110001100100011000001010001111011001111110010011011111111111101110001111001000100001110000010011111101110010000111100000111011001011110010100101110101000100001110010010001010100111111011111000010010010111111110001100111011011011000010110101100111010010011010100000001001101000011101000100010110001100110101110000000011110000010110110111010001111100100001110010111001111101011010100010010111100001010111011101110110000101000000000011100000000100110000100001010110100111111001011010111110101010001001010001111111110001101011100110000010001010000101011111110010000000100000110100100011110011110011111000110011000000000011001110011000000000110111000001011111110101101000101000001111000101110111110001111110011011011010100000000100000100011111010001100001001110000110010000110100010010001000110011000000111111111110011111100010000111111100011010100111001111100001010001101011011100000100000011010111000111011101011110111010010000101000011000110111001001010000101001110110011101001000011010110011001111110101000100001110001111100000101100011011001001000011111101100111100101011111100110110111111000000011010110011010011000000100010110110110011110001110101100100111001011110110000100000101100000111100111101001011111001111111011101111100001100001100111001000000110111100111100011101001111001010111111010011110110001110000000000010001111000011100100111100110100001001110010011101011001011001010001101101101110111011001000100111000001111101001111000000110110100101110001111111001101101111111000110010000100010110010011011111001101110011100111100110001010100111110110010001100011111001101010011011000011111111111001001011100010000001000110101011000000101000111011100100011000100101000110101100001000011000000010010110001101101001101010111100111001001111111000111101111000100000000001111101110011101001000010111111000000101011001111110011000000100011101101011100011111111110010000000100000100011000100001110001000001000110100110100111100111101010011000001001111001101101000111100000000111101101000011110101100000001110100001100001101001101001001111000100111100000000000111100001110111110111001111011001100011001011111010000111101110010100001001101101110101110000100100011000110010111001000011011111011100101110110100001000100011100100111000110000000101000001110110000101101100100000100101110001000011010000110001000101001010011100001101101010001111101101000000111110011101000110101001000100011000001110111111010001110100100110110101111111101111000101111110100011101111100000011001100111000000110001111111100010011100101101110110101010000101001110111011110110110100111110110001110111101100001100110000011111111011110010111011011100000011000101001100110110110100110010001010010000100010100011101100000001011010111110010111010010011101000111011110010011111000111011110000110100101100111000010010100000101001001011010101100010011011101011010111100110011110100011000110000011111101110000110011100000101011001011101000011111001111000010000100010111001001001111011101110000011100101001011100100010101100000111011110100111100101110000101001001110101101010001111001001100010001110000101100101101110000000011001100000110101100111011011011010110110001110110110011001101101100101000000010000010101001000110111110100110011111011100100110100011100001101110000001000101100010011101100011110000001010110111001110110011000100111010010011010101110000001111111011101110001001110000110001011100001100110001101111011010001100110100001001010111111000011101111111100010001011000010001111000111001011001111101111000010011100000000010001011111110010010111101000011010110001000110100011011111110010111011110001100101110001001110011110100100111011110000011011000000000010010110101101000111100101000111111110000000011100100100101010110000001101010111001100010001110011111111001000001010111111010100100111000000111010100001001110111011010010011010000000001011111100111010100110001100010100101000001000000110110110001001010001101100000111010100011001111011101111100000110100100110110101010001000010110100000011000000111100000000001001010110011010101100101110101011111001110000110001111111110001000111111010001101100010001010011000001011000000110000100110111111000001101100111110100011111010110111101101000100000001010111011100011101111100111000101111100110110000001000010011010100111000010011110100111100111000111100001111101000000001011100010000010100010011000001001010110011111000000100100101111111011011111100000000110111000000100111000000000110101101111101010001111000000100100111011010001000010000010101111111100011101111101101100000111011001010010000111011010100111100000010110011101110000000000101000111101010101010001100001001011001011100000000001001000001110010001000101101101110001010001011001111000101001001010100111110100000101001100111111011100110001000000001000110000001100000011001110011111101100110100001000111001110111111111101100011110111000000001101111000111000001101000001110111110010101101011101000100110011000111100110001101000001011011100011010101010000010100110010001110010010110000010001000110011001110001101011111011110010010010000001110111000010000000111100111101101001010000001100000010000001111101001111001101011110011000011011111111100001000000001111110110001101010100110111000101110;
localparam PROTOTYPE_LEFT = 10000'b0111000101111000011110111100111111100001000001111111000110111100101111110100001011100010100000111100000000011010111010110010100011011111010000011100000110001111000111100010100001110100000110010111010101100101011110101100010000101000111101101110001110010001110011110000111110001110010011001000100000100001100000000100110110100000100000001100011100000110001110010010011000111110011011100000100100100110101100111001001101000000110000010000000011000100110001101101001100100000011101011011100010011101110010111111111000100000000111100100100011001111010010111110100010010000101000001101110011000000100111011000101101010001101011111111101001100101111110001101011111110111100000100011010101100001000011000001000100111110100100110010111111101110110011000001111100101111110011111110000111011111011101110110000100000111100011001000111111001101111111100100110000100100110011001110000001010011001111100111001111101111000111101001100111001100010111010011000011000111111111101111110110001000001011010110101100100010101001011111110011111010110000000011101101111011000000101000110010110000111101110011000011110111111000011111110100010000011000011101000110111000101010011000011100011110100110111011110001010000110111100100000110100110001000111001010101011101110010111100001110000001100001000001110001000011001100100000000100011100000111011010001000011101110001011011111011111111101100101000111010101011010010100111100101111000101010000001011111111111110011000111111001100100111101001000100001101101001011000111000010100010111110011111101000111011011101100000010010101000011000101001111101100111011100010111100100000111000011011011111000101100011000011111011101000100100101001111000000100100011111111110111110010111011110001110010101011111101001100011001111000000111110011111110100000110001001111110100101110001010001110110011100001000000111110011100110001101101100111010101101111011011110001101001111100111111001100011101111111110010000101111001111100111011000000100001111011110110011110101101101011011110001100001110111100000111100010111101010100110101100001010001101011010101101101111110100010001010110101101000010001010000111000000010011001011110001011001100101100001101101110000011011111000000011000100100000011111010011000110110000000001111011100110001100000010011110100111010111011101110110110110110101010011111110010110101000101010110011000110110110011110000101011001100000001110101000011110000010100111100011110011110000111110101001110011100000100001001011010101100100100001000000011000100110010000001101100111100110010010000011101111011110111010100010000011111001000111011000011101100010101110101100110000011100001010001010000001100001001111101011110110010001011111101000010010010000111011011100111000111011111000010010110001010111010001111100111110110100000000001001111100000111010111010110111110010111000000011110111101001011000110010011000011110000101010111010011111100000000101011001010000010100011011101000010010010111100101011101010100101111111000110011110101100110110111001100010111100110001111000011001100100000100011001011110100101001100111010010110000000001101100001010010000100010011100111111010100110111100001010001010001001000111111110100000000100010100100001111011000101101111011110110001000101110000000101100110010001111000001101010110011101101011000111110001000010101001101110011110001000101110100011011100010011001000111111001010111100101101110011101000100111111011100010010100010001110001000110011101111011100111111101101100100001010001000011001010000011110001111111000001101011100000001011111001110100111011011000010100010101000100010101100001110001011110000001111011100111001010100010011101010110100000011011010011110000011111000110001100011001100111101011001100101000101001011000000011100011000111110000101011100010000001000000111011001011010000010110011011111011000000100000111111011011000101001011000001100111110000000111000110111101111101000110010100100000111110011111010101011011001000010011011000100001110001001001100000011111111010010010100000000010000101101011101010110100111101111010001000001100010011001011000001010100101101101111101010001001101010000110111010100000010100111010101000111000001010000001111110110101011110110100000000000111011101000000111001011010001101000110001111100010011111101010011100101001011001110010100101011000111010100100010101101111000010010110100000110001001101010110010011101110001011111111111011001100111100001110101101010000000110111000010100000011101110100111101110111110000111001100000100001110000111011011011000010000001100100000000111111000001000001101000101010111101110101101010000000000110011010100110100000010100010110000011001011101000011100001100000001000111111111101111000111010011110001111100101010000011011101111000011011100101111011011001010001000110101011001011111100011110010001000001110010011111110001010000100101001000001010000111000100001111001111110101010011111100100101111000001010001111011000000001010011000111111011101110001111001111000001100000010011111101110010000011100010110011000011100010000101110101010101001110010011011010100111111011111000010010010111111000101100111000010101000010001101100111010011100010100100001001101001100011000100010110001100001101110000000001110000011001110111000011111100110001001110111001010010001010100010010111100001011000101101110111111101000100000011101110010101110111010100000110100110111000100010111110101010010110010001111111110001101001100110000010001011100101011111110010000000000001110100100011110011110011111000001011000000000011001111110000000000110110000001111111110101101000001000000111000010110111110001101110100100110000001000000100100100011010001001100001111110000110100011001100010010001000111010111010111111111011011111100010111111111100011010100111001101011111101111101011011001111000001111110111000001011101000010100000010000001000011000001000001110111000101011000100110100110110011010110011001111110100000111001110001111100001000100111111001001100011111110001111100101000001100110110110011111100011010111011010011000000100010110110110011111111110101100101001001011110100000100000101000000111100111011011011110001101100000010011010111100001101000001100000110111100101100011101011011010011001111011111110000001111011000000010001111111000110011111100110101011001110010011011001001011011010111101100011110101011001000100111000001100001001111111110110110100101110001111101001101101110101000110010000100010100101000011101001101110011100111100110011001101001110110010001100111111000001010011101000011111001011001101011100010000001001110101011000000100000111011100100001011001001001110100100011000001000001011001001111101001000100101111000111001001111111000111001111000101010010001111101110000101011000010111111100000101010001111110011000000100001101101011100011111111110011000000000011000010000100001110001110001000100100110100101101001101010011000001001011001101101000111001000001101001100000000110101000111000110000001101111101001101001101110110100000100100000010101101000001000001111000000010111100011001000111001100111101110010100111001101101110111001010001100001000110010111001100011011111011100101110110100011011010011100000111001100000000101000001110100000000011111100000100011010001000011010000110001010101001010011100001101101010001111101101001100111110011001000110101001110000011111001110111111001111100100100110110011111100011111000100010110000111101100111000000011100111001000110000011000100010011110101100010110101010010110001110111111101110110100111110111101110111101100011100000001111000111100000010101010011100000011000100001100110001110110110010001010110000100011100011101100000001011010111010001001100010010110000000111101010010111000111011110000110101101100111000000110100000101001110011010111100010011011101010110001010001111110101011001110000011111011110000110011101000101011001011101001000111001111100010000100010111001001011000011101101001111100011001111100100011101100000111011110100111100101110000010101001111011101110001110111001000010001110101100100101101101110000011101100000111000010111100011011010110100001110110110011001100001100100000000011101010101001000010101000100110010011000100100110100011100001011110000001001001001101011101100100010000000001110100010010110011001000111110010011010111110000001111111111101110010001101100110110011100001100101001101111010100001100101101001001110111111100011101101111110110101011000011001111000000001011001111101111000010011100000010010001011111110001110101101000011000111001000111100011010000010010111011110001111001110001001110111110100100011011001111010011000000100010000110101101000111100110000111111110000000011111011100100001000000001101010111000100110001110011110111011010100010111111011100100101000001110010100001001111000100010010011011000000001001111100110010010011001100001011101100001010000110110110011011010001101100110111010100011001111011101111010000110100100110110101010001010010110100000011000000111110100000001011100010011010101100000110010001111000100000110001111100100001010111111010001101100010011001001000001011011000100000100110111111000001100100001001100000111011110111101100000100110001010111011110010101111100111000101100000000110000001000110111110101000000010000111100111100001110111100101000001000000001000011110000010000010011111001000010010011110110111100100101111111011011101100010000110001011011001111000010000110101101111101101101111000000100100111011010001000010000011100001111101010001110001101100100111011001010010000111110001100111000000010110011101110000000100101000111101000101001000010001001000101011000101000001001000001110011011100001101111100100110001011101100000101001001010010001110000000000110000111111011100110001000000001000001101110011110011100001010011101100110111001000111100110011110101100100011110111010000010001111000111001001111000001110001111010001101011101000000100011000101110110001101000001011011100011000100010100000011000011111110010110110000001101011110011001101001100011111011110010010011000111110111000010000000111100110101101001101000001100000010000010000100001111001101011110010011011000101100000001000000001111110110011111000100110111000101110;
localparam PROTOTYPE_RIGHT = 10000'b0110000111111000011110110000111111100001000001111111000110111100101111110100001011100011010001011100110001111000111010110010100011011110010000011100000110001111000111100010100010110110000110010111010101110101011111101100010000011000111101111110001110010011110011110000111110001010010111001000100000100001100000000100110110100011000000001100111100000110000100110010111100110010011011100000100100110110101100111001001101000001010000010011000010000100110001101101001101101000011101011011100010011010110011101111111000100000001111110100100010101111010010111110100010010000101000001101110011000100100111000110011110011001101011111111101001000101111110001101011001100111100011100001010101100101000001000101000100110010101011110111000011101110010011000001011100101111110011111110001111011111011101110110000100000111100011000000111111001101111111100100110100100100110011001110000001110011101111100111001111111111000111101001100111011010010111000011000011000111100111101111110110001100000011010100101100100100101001001111000011111110110000000001101101111011000000101100110010110000111101110011000011110111111000011111110100010000011000011101000110111000111010011100011101001111100110111111110001010000110111111100000110100100010000111001010101000001111101000100001111000001100001000001110001000011001100100000000101011111000110011010001000011111110001011011111111011111101100101001011001101101000010100100100101111100101010000010011111110111110010000111111001100100111101001000101111101011001011000110000010100010111110010110011000111011011111100110010010101000111000101001111101100111011100010111100100000110000011010110001000101100011000011111011101110100100101001111100000000000011111111110111110010100111100001111110101011111101001100011001111000000111110011111110100000010001001111110100101110001010001110110011100001000010111110011100110110111110100111010101101111011011111101101001111101011111001100011101111111110010100101111001111100111001000000010000111011110110000000110101101011111110001100101101011100000111100110111101010110111000100000010001101011010101101001110110100010001010110101101000010001000100000000000010011001001110001011001000101110000101101110000100100001000000011000100100000011111010011000110110000000010111011100010001100000000000100100011010111011101110110110110110101010000111110010010101000100010101011001110100110001000000100011001100000001111101000011110000000100111100011110011110000111110101001110011100000111011001011010101100100100001000000011000100110110111110101100111100110010000000011111111011110101010100010000011011001000101000101011111100010001110101100110000011100001010001100000001000011000011101011110110010001011111101000010010010000111011011100111011111011111000010010000001010111010001111100011110110111000000001001111111000111010111010110110110010111000000011110111101001011000111110011000000000000101010111010011111100000010001011111010000010100011011101001000000010111100101011100001100101111111000110011110101100110110111001100010111100110001111000011101100100000100000001011110100101001100001010010111000000001101100001010010000100010011100111111011100110111100001110001010000001000111111110100000000100011100100001101011000001101111011110110111000101110000000001100110110001111000001101010110011101101000000111110001000010101001111111000010001000101110100011011100010011001000111111001010111111111001110010101000100100010000011010001100011001110011000101011111111001100100001101101100100001010001000011001010011100001001111111000001101011100000001011100001010100111011010000010100010100000100010100100011110001011110000001111011100111001010100010011101010110100000011011010011110000011011000111110000111001100111101011101100101000101111011000000011100011000111110000101010101010000001000000101011001011011000010110011011111011010000100000111111011000000010001001000001100111110101100101101110111101111101000110010100100000111110011111010001011010111000010011011000100000110001001001100000010011101000101110100000000010000101101001001010110100011001111110001000001100010001110010000000010100101100101111101110001101100011110010101000110100010100111010101000011000001010000001111110111101111110110111100000000111011111000000111101011010001101000110001111100010111111011010011111101001011000110011100111011000111010100100100101101111000010010110100000111001111000110010010011101110001011111111111011001100110100011110001011000000000111111000010100000011111110100111101110111110000111001100000100001110000001011011011000010000001100100000000111111000001000010100000101010111101110101011010000000000110011010100010100100010101010010000010001010101110011100001101100000111011111111101111000111010011110001111100101010000011011101011000011011100100111011011001010001100110101011001011110100011110010001000001110011100111110001010000100101001000001100000111000000001111001111110101010011111101100101101000011010000011011000000001100011000111111011101110001111001110100001100000010011111101110010000011100010110011000001110010000101110101010111001110010011011010100111111011111000010010010111111001111100111000111101011010001101100111010010100010100100001001101001100011000101010110001100110101110000000001110000011001110111000011100100110001001110110011010010001010100010000111100001011000101101110001101101110100000011101101010101110111100100010110100110111001111010111110101010010101010001111111100001101011100110000010001011100101011111110010000000100001111100100011110011110011111000001011000000000011101111111000000000110110000001011111110101101000001000000111000010100100000000101110100100100000101010000100000100010111010001100001111100000110100000001100010010001000110011001010111111111011011111100010111100011101011010100111001101011111101111101011010101111000000011110111000110011101000010101110010010101000011000101101001110110000101011010100110100110110011010110011001111110100100101001110001111100001000100111111001001100011111110100111100101000001100110110110011111100011010110010010011000000100010110110110011111101110101100100001011011110100000100000101000000011100111011011011110001101100000010011011101100001101000001110000110111100101100011101011001010011011111011111110000001111111000000010001110111011110100111100110101011001110010111101011001011011010111101100011110111011001000100111000001100001001110111110110110100101110001001111001110101111100100110010000100010110101000011111001101110011100111110110010101101001110110010001100111100000001010001001000011111111111111101010100010000001011110101001000000101000111011100100011011001001000100110100101000010101101010101001111101101000010100111000111001001111111000111101001000100100010001111101110011101011000010111111000000101010101111110111100000100010101101011100011111111110011000000100001000011000100001010001111101000100100110100101101001101010011000001000011001101101000111101000000111101101000011110101000110000110000001101111101001101000001111010100011100100000010101111000001000001111110000110111100011001000111101100100001110010010110010101101110111001000001000001010110010111001000011011111011100101110110100111010100011101000111001110000000101000001110110000000001111100000110011010001000011010000110001010101010110011100001101101010001111101101001100111110011010000110101001111000011111001110111111001010000100100010110101111100011111000100010110010111101100111000000011100111000000110000000000100010011000101101110110101010010110001110111101101110110100111110111001010111100100011100001000011000101100000010111011011100000011000100001100110001111110110010000010110000100011100011101100000001010110011010000111000010010110000100000001010010111110111011110000110100101110111000000110110000101111001011010011100010011011101010110001010001111111010011011110000011101101110000110011101000101011001010001000001111001111000010000100010111001001011000011101101001111100111001111100000000101100000111011110100111100101110000010101001111011001110001111111001000010001110101101100101101101010000011001100100111000110111100011011010110100001110110111111001100001100101000000110010010101000011010101000100110010011000000100110111111100001011110000001101001101111011100100100010100000001110011010110110011001000111110010011010101110000101111111111101110000001101100110110011100001100101001101111010100001100101101001001110111110100001101111111111110010111000011101111000000001011001111101111000010011100000010010001011001110010010101101000001000111001000110100011010000010110111011110001111001110001001110111110100011011011001111010011000000000010000110101101000111100110000111111110000000011111011100100001000000001101010111000000010001110011111111011010000010111111010100100111000001110010100001001111010100110010000010000000001001111100110010000010001100010101101100011001000110110110011001010001101100011101010100011001111011101111100010100100100110110101010001010010110100000011000000111100100000001011100010011010101100101110110001111000100000110001111111100001000111111010001101100010000101001000001011000000000001100110100101000001100111101111100000111011110111101101000100110001010111011110011101111101000111101100000001110000001000110111110000111000010011111100111100111000111100001000001000000001000011110000011101010011111001000010000011111110111100100101111111011011101100010000110011011011001111000000000110101101111101110101111000011100000111011010001000010000011101001111101010001100011111100101101111000000010000111010001100110010000010110011101110000000100101000111101000101001000010001001001101011000001000001001000001110011011100010010111110011010001011100100000101001001010010110000100011101100000111111011100110001000000001000001101110011110011000001011111101100110111001000111011110011110101100100011110111010000001001111000111000001111000001110001111010001101011101000000110011000001100110001101000001011011100101010111010100010100110011111110010110110000000001011001111001101001100011111011110010010011000000010111000010000011111100110101000000101000001100000010000010011101001111001101011110011000001000101000000001000000001111110010001101010101100111000101110;
localparam PROTOTYPE_YES = 10000'b0111000111001100010010110000111111100001110001111111000110111100101101010100101011110011010001011100001001011001001000101011100011011110110000010010001000001100001111100010100010110110000000101000010110011100011110101100010000101001101101101110001110010011010011110000111100001010011100001000100000100001101100000100111110111100110101001100011100001111101110010010011000110010011011100000100100110110101100111001101101000001010000010000000000100100001001101101001100100011011101011011100010011101110001111111000110001000100111101000100100101101010010111110000010010001001000001101110011000000111100111000110011011001100011110111101011100101111110001100010111100111100011100011010101111110001000101100100100111100000011110001000111100010001100010111001100101100110011111110011111011010011101110110000100000111100010100000111111011101111111100100111100100100110011100010000001010000101000000001001111100011000010000011100111001100010100001111000011000111111011101111110110001000001010010100001101100000101001010001110011111110111100011111100000111011000000101100110010110000111101110011000011110111111000011111110101010000000000011101001110111000101010011010010000011110011000111111110001000001110101111100000110110100010000111001000111011111110010111100010000000001100001010001110001010011001111111000010101011111000000101110001001111101110101011011111011111111101100101001011001111011010010100000001101100100101110000001010111000111110011000111111001100100111101001000100001100100001011000110000010100010111101110001100010111011001101100011010010111000011000101001111101100111011100010111100101110100000011110010111000101100010000010010011101000011000101001111011000100001011111111110000000010110011101101111100101001011001011100011001111001000111100011111110100000000001001111110100101110000010001110110011100000100011111110011111110110110101100110100101101010011011100001101001111100111111001100011101111111110010000101111111011100111011000000100001111011110101111110101101101011011110001100000110011110000111100110101101010100110110100110010001101011010101101011110110100011111110010101101000010001010000110000000010011100001110001001001000101100100101101110100010000101000010011011010000000011100010011000110110000001001001011100010010100010000001110100011010111011101110110110110110111010011110110001101101000110111000111111010000010001001101100011001100000001101101000011010000000100100000011110011110000111100001001110001100000100001001011010110000100100001000000011000100110010111111101111011001110010000001000101110011110010010100010000111111111110101001000011111100011110100101100111000011000011110000010000001100001001111101011110110010001011111101000010010010100111011011100111011111011111000010110110001000111010001111100000010110111100000000001111100000111010111000110111110010011000000011110111110001010000110010111000111001000101010001010101111100001111011000001010000000100111011100101000010100111100101011101001100101111111000100011001110001110110111001100010101100110001101000011101000010001110000010011010100101001100001010010110000000000100100001110100000110010011100111111010100110111101100110011010001101000101110111010000000100010110011001001011000001101111011110110111110111110010001001100110111101111000001101010010011101101011000111010111000101010001101110010010001000101110110011011100010011001000110111101010110000010101110011001000101100011011111010011100011001011100010101011101110010100111111101101100100001010001001011001010000011110001111111000001101010010000000000011001110100001111011000100100010111000100010100100001010000011110000001111001100101001010100010011001000111100000011011010111110000011111000111110011011000100111101000101100101000110100011100000011100001000111110000101011110010010001000100101011001111011000000100011011111011000000100110111100111011000001100111000001100111110100000110000110001101111101000110010100100000111110011110010001011001000100010011011010100000110001001001100000010001111000101010100010000010110111001001000000110100100101110110001010001100010011001011001000011001001111001111101010000001101010010110101100100100010010000110111100011000000010010000111111111101111110110111111100010111011111000000001101000100011000000110000010100010010111001110001111100001011001000100100101010110001010100101000110001011000010010110100010111001011001110010010011101110001011111111111011001100111101011110101001010000100100111000010100000011101110100111101110111010000111001100010110001110001001011011011011010000010100110000001000110110011000001001001001010111101110101011001000000000111000000100101100110111101010011000011001010011110010101001100000000111001111111101111010100110011110000111100101010001111011101010000010111100101111011010001000001010110100101001011110100011110000001000001110000101100110001010000100100101001001100000101000000001110001111110111100011100101100100011011011010000011011000100000010001000111111011101010001111001110011001100000010011111100110010000001101110111011010011000010100100110101010101000110010011001010100111111011111000001100000111111100011100111000110100111010001101101111010011100010100100001001101001100001000111011010001100110101110000000001110000011111110111000011101100110001111000111001000011010010100010010111100000001000101101110001111101001000010011100000010101100111011100011110100101111010100011111110001010010111010001111111110001101011100001101101001011100101011011110010000000100111111100100011110011110011111000110011000000011111101110010000000000110110100001111111110101101001110000001111000101000111111111001110000100100000101000000000100100001111010111000001110001100000110100100000010010001000111010110010110011111110011111100010001100011101001010100111001100111001110111101011010000110000001011110110111110011101011110111100010010101000011000001000000110111000101011100110011100000100011010110011001111100001100000000110001111100001010000101110000101100011101110100000000101011111100110110110011111100011010111101010010000000001110110110110011111101110101100101001001011110101010100010111111110011100111101011011011101101100000010011010101100001101000001100010110111100111100011101001111010011000001010011000110001100111110000010001110001111101100111100110101001001110010011101011001011001010111101100011110110101001100100111000001111001001110110000110111011000111011011111010110101101111000110010000110010110100000011110000101010011100111100110011000100111010110010001100111101000011011011101000011111001111000001010001101100001001000101011000000100000111011100100011001010001001100100100101000110101101011101101111101101000001000111000111001001111111111111101111000100010010001111101110011101011000010110111110000101011000011110010000000100000101101011100011111111110011000000101100111100101101001101001111100000110100110100111100001111000011000000101110001111101000111001000101000001100000011110101000110000001000001100000001001101001001111001100111100000000000001110000001000000101110000010111100011001000111010100000111110010000011001101101110111111010111100001000110010111001000011011111011100011110110110001101100011100000111011001011110101111101110000000000000011110010100010111001000011010000110001010111010110011100001101101010001111101001001100111110011101000110001001000000011111001110111111010000000100100100110101111100011111000100011110000101010010110000000011100111001000110001111100000100011010101101111110101010000101001110111111110110110100001110111000010011111100101100110001111000111100000010101011011100000011000100001100110110110110110010001011001100100010100101101100000001010100011011100100111110000110001000101101010010111100111011110000110100101100111000010110100000101001001011010111010110011011101011010001010001111110110011001110000011111011110000011100011000101011001011101000001111001111000010000100110001000111101001011100101110000101111001100000001001101100000111011111100111100101110000100001001110111101111001111110001100010000000101100100101101101000000011001100100111000110111100011011000110100001000110110111001100001000110000001000000110101000000010000110000101111111011000100110100011100001011110000001001001001100110101100011110100000001110010001010110011000000111110010011011100110000001111111111001100011111101110110111000100001000100000101111100000001110111011000001010100010100011101111111111101010111000011001111000000000011010001101001101100011100000010010001011111110000110111101000011010110001000110100011010100010010111011100001111001110001001110111110101111011011001111010011000000000010010110101101000011100110101111111111000000010111011100100001000000100101010111000000010111110011110111011010100100111111001000100101001001111010100001001000000100010010011010000000010011111101010011010111001101001100111100001001000110110110011001010001100100011111000011111001111011011111011001100100100110110101010001010010110100001100100010101010100000110010000110011010101101101000001001111000100000110001111111100001010111011000111101100000001101001000001011000000001100100111011111000001100111111101000000111011111111011110111000000001010111011110111101111100111000101100000110100000001000000011110011000100010000111100111100111110111100001000101000000001000011110000011100110011111001000010100011111000000100101001011111001010100000000000110011101000100111000000011001101110111101101101111000000100100111011010011101110011011100001111100001001111101101100101111011000100010000111011100100111000000010110011101110000000100101000111100111001001001100001001001101011111101000001001000001010011011100010001110001000110001011000100000101001100010101001110100010110101111010111011100110001000000001000001100110011000011100001011111111111010011001011111100110111110111100000011110011010000000101111000111001110110001001010111111010001101011101000110110011000101100110001101000001011011111101010011010100010100110010001110010110110000100001011010011001101101100011111011111100010010000001110011000010000100111100110101101100100000001100000010000010010011001111001101011110010000100011101000000001000010001111010010011111010011000111000101110;
localparam PROTOTYPE_NO = 10000'b0110000110001000010001010000100000100001111001111111100100111100101100010100000011101011010000111100000001011010111010110101110011011110010000011010000000001111000111100010100010110110000110010011110011111101001111101100010000101000111101001110001100010001110001110000111110001110010011101000000000000001101100001100110111000011000000101100011101111111101110000010011101011110011011100000100100110110011100111001001101000000100000010000000010011110110001101101001100101011000101111011100010011001110010111111001000000000100111110110011011001110100010111110001101110010101000001101110011000001100100101001010010011010011010011111100010100101111010001111010111110111100011000011000001100001000000000100100100111110101011010000111100100110011100100001011100101111110011111110000011011111011101110110000100000111101010001000111111110101111110110101110100100101110011000110000001010011101011100111001111100011100000010111100111001100001000100011011101000111111011101111110110001001000010101000111101100000101001000001110011111010110011100001101111111011000000101100110010110000111101110011000011110111111000011111110101100100111000011101000110111001101010001100110000011111101110111111110001000001110101100000011010100000001000111001011101000111110010111101101111000001100010111110010001000011001111111110010101000000000111011110001000011111110001011011111011011111101100101001011001101011110010110000010101111100101010000001011111000111110011000111111001100100111101001000101111101100001011101110000010100010111110011001101000110011000100010110000010111101111000101001111101100111011010101011100100000100000011010110000111001100011000011111011101000100100101001111011000100110011111111110101111010111011110011110010111011111111110000100001111000000111110011111110100000111101000111110100101110001010101110110011100000110000011110011100001110111101100110110100001000100011100001101001111100111111001100000101111111110010100100111111111100000010000001000000111011110110010000110101101011100111110001100101010010001100100110101101010100111000100110010001101011010101101011110110100010001010110101101000111001010000000000000010011111011110011011001100010100000101101010000011011110110000001000100101000000100110000000110000000001001111011100110001100000000110010111011000000011101111110110010110101010011001110010011101000101010110011000110110110001110110101111001100000000101000000011110000000100111100011110011110000111111001001110011100000111111001011010110000100100001000000101000100000010000001101011100000110111010001011000111011110010010100010000011111001000100111010011101100011101110101100110000011011101010001000000001100001001111101011100110010001011111101000110010010010100011111100011001100111111111101110110010110011010001110000111110110011101100000001111100000111010000100111111110010011000000011111000101001011000000010111000111111000101010000001101111100010011010000001010001000100111011101000001110010111100101011100001100110111111011010011110101110110110101001100010111100110001101000011001111100000100111101111110111011001100001110010110000000001101100010010010001110010011100111111011101010101110001001101010000001100101110111000000001000111110100001110011011101010000111010110001101100110000010101100110110001111000001101010010011101101000000110101001000010101001101100111110001000101010110011011100010011001000111111000100101100101110000011101000100100011011111010010100011001110100110101011110011010100100001100001100100010010001001011110010000011001001111111000001101010000000000100001010000100001010011000010100010101000000010111100001110001011110000001111011100101001010100110011001000010100000011011110011110000011111001001000100101001100100001111100011010110101101011000000000000011000111111100101000000010000101010000100011001111010000001000011111111011001000111000111111001000001101010010000000000111110000010110000110111101111111000110010010100000111110011111011011011001111010001010000100101111010001000001100000011000111000101001100110110010110110001001000001001111100111101110001010001100010011001011000001011011101111010111101110001001000010100110010110101000011111000110111100011000001010000011111110010101111110110111111100000111010001000000111101000111100000000110010111100010010111101010011111101001011001110011100100111000111010100100000101101111000010010110100000111000001101010110010011100011111011110000111011010110111100000110001011000000000110111000010100000011001110100111101110111111111000001100001000001110010111010011011100110011100100110000000111111000000010001101011001010111101110101010011000000000110011010100100100100000100000110000011001010011110011100001101100000111011111111101100101000010000010001001100100011000011011101011100100111100000111011010001101110110110100011111011111100011110000001000001110000011011111001010000100101001101001100000111000000010010011001110101100000110011100100011000001010001011011000001000010011000111111111101110001111001000100001100000010011111101110010000101100000111000001011110010100101111011000100001110010010011010100111111011111000010010010111111110001100111000011011000010110101100111010010100010100100001001101000011101000100010110001100000101110000000011110000010111110111010001111100100001110010111001111101101001010010010111100001010111001101110110000101001000000011101000000101110000100001001110111110111001011010111110101010001001010001111111110001101101100110000010001010000101011111110010000100000000110100100011110011110011111000110011000000000011001110011000000000100110000000111111110101101110001000000111000101110111110001101110011011011111100000000100000100011011010001100101111110001111011000101100010010001000110011000000111111111011011111100010000111111100010010100111001111100111011011101000011100000100000111000110100110011101000010111010010000001000011000110111001001110000101011101110011101001000011010110011001111110101000100001110001111100000101100010011001001000010111101100111100101011111100110110111011100000001010111011110011100000100010110110110011110001110101100100111001011110110000100000101000001111100111101011011110001101111011101111100001100001100111000001000110111011111100011101011011010010111111010011110110001100000110000010001111111000110011010011110100001001110010011101011001011011010011101101101110101011001010100011000001111101001111000000110110100101110000111111001001101111111000110010000100010111010011011111011101110011100111100110001010100111110110010001100011111001101010011011000011111111011001001011100010000001000110101011000000101000111011100100011000101101000110101100011000011010010011010101111101101001100010111100110001001111111000111101111000100100000001111101110011101001000010111111110100101011001111110011000000100011101101011100011111111110011000000100000100011000100110110001000011000110100110100111100111101010011000001001111001101101000111100000000111101100000100110101100100010110100001100001101001101001111111000100111101000000010001100111110111110101001111011001100011001001111010000110101110010100101001101101110101110000000100011000110010111001000011011111011100101110110100001011010001100100011000110000000101000011110100011000101100100100001110010001000011010000110001000101001010011100001101101010001111001100010011000011011011000110101001000100011000001110111111010001110101100100110011111111101111000101111110100111101111100000011100000111001000110000011000100010011110101101110110101010000101001110111011110110110100111110111010010000101100001100110000011111111011110010101111011100000011000100001100110110110100110110011010010000100010100011101100000001011010111111100111010010001101000111011110110011111000111011110000110100111100111000010010100000101001001011010101000010011011101011010111110001011110101011000110000011111101110000001011100000101011011011101001000111001001011010000100010111001001001001011101110000011100101001011100100011101100000111011110100111100101110000101001001110111101000001111011001000010001110000101100101101100000000011001100000110101000111011011011011010110001110110111011001101101100100000000001101011101001000010111110100110011111011100100110100011100111101110000001000101101110011001100011110000001001110101011000110011000100111000010011010111100000001111111011101110001001110000110011011100001100100001001111011010001100110100001001010111111100111101101011100011001011000010001111110111001011001111101111000010011000011100010001011111110010010111101000011010110001000111100011011111110010111011110101100101110001001110011110100000111011110000111011000000000010010110101101000110100101000111111110000000011110000100101110110000001101010111010100000001110011111111011000000010111111010101100111000001111010100001001110100011010010011010000000001111101100111010100011001000010100101000001110000110110110001001011111101100111111010100011001111011101111100000110100100110110101010001000010110100000011000100111110000000001001000110010010101100101110101011111000000000110101111011110001000111111010001101100000001010001000001011000000110000100110111111000010101100111110100011111011110111101101000100000001010111011100011101111100111000101011011000110000001100000011110100111000010011100100111100111000111100001111101000000011111100010000010100010011111001000010110011111000000100111001111111011011101100000000110111000000100111000010000110101101111101010001111000000100100111011010001000010000000101101111101000001011101101100000111011001010010000111011101110111100000010110011101110000001000101000111101010101011001101011001011001011000000000001001000001110010001000001100111110001110001011001100000101001001010011011110100100101001100111111011100110001000000001000110000001100000011101110011111001100110111000000111101110011111111101100011110111000000001101111000111000000111000001110111111010101101011101000110110011000111100110001101000001011011100011110010010010110100110010001110010010110000010001000110011001110001100111111011111100010011000001110111000010000000111100111101001001010000001100000010000001111101001111001101011110011000111011001111100000000000001111100010001111110100010111001101110;
localparam PROTOTYPE_UP = 10000'b0110000011111000011110111100111111100001000001111111000100110100111111110100001011100011010000111100010010011010111010110101110011011111010000011100000110001111000111100010101101110110000110010111010101110111010001101101101101010000101101111110001110010001110001110000111110001100010011111000000000100001100000000100110101100011100000001100111100000000001001100010011101010010101011100000100111100110011100100001001101000000100000011000111110000100110001101101001100101000010101111011100010011000011010110111111000100000001111110100110011001111010001111110000010010000101000001101110011001000100111101000010000010001101011111111101001000101111110001101010001100111100011100001010001100001000011001001000100111110101011110010111100101111110011000001011100101111110011111110000111001111011101110110000100000111101001001000111111001101001110110111110100000000110011001110000001110011001111100111001111101111000101011011100111001100110011100011011101000111000111110111110110001101000010101100111101011110101001101110000011111001110011100001101101111011000000101100110010110000110101110011000010000111111000011111110100010000111000011101000110111000101010011100010001010110000110111011110001011100110111100000000110100100001111000001010011011101110010111101101111000001100001000001110001000011000000000000000100011100000111011110001000011111110001011011111011011111101100101010111010100111000010010000010101111000101110000000011111111001110010000111111001100100111101001000001111110011001011001111000010000010111110011110011001111011011111100110010010111111111000101001110001100111011100010111100100000111100111011011101000101100110000011110011101000100100101001111011000100110011111111110001110010111011110001111110101011111100001100011001111000000111110000111110100000000001001111110100101110001010101110110011100001000000011110011100110001101101100111010101101111011011111101101001111101011111001110011101111111110010100101111111011100111011000000010000111011110110000000110101101011100100001101111001110000000111100010101101010100110111100001010111101011010110011101111110100010001010110101101000111001001000001100000010011011001111001011001101010100001101001110000011011111000100011000100100000011111010010000110110000000010000011100110001100000000111010111011001000011111010110110110110101010011001110010010101000101010110011011110110110001110001110011000100000000111100000111110000110100111100011110011110000111110101001110011100000111011011011110101100100100001000000101000100000010111110101100111100100111011000011011111011111101010100010000011111001000100011010011101100000001110101100110000011100001010000110000001100011001111101011010110010001011111101000010010010000111011111100001001111011111000010010000001010111010001111100111110110100000000001001111111100111010111010110100110010111000000011110111101001011000000000011000111001000101010111010011111100000000010100101010000010111011011101000000010010111100101011101001100101111001011110011110101100101100111111000010111010110001111000011001110000000100111101011110111011001100111010001101100000001101100001010010000100010111100100111100101010111110001001101010000001111001110111000000000100011100100001110011011100100000111110110111000101110000010111110001010001111000111101010110100001101011000111110001000010101001011010000010000000101110100011011100010011001000111111001000111100111010000010101001000111011011100010010100010001110000010110001010011001100100001101101100100010010001001011001010001000001101111111000001101010010000000100001001000100111010010000010100010101000100010100100001110001011110000001111011100111001010100010011101010110100000011011010011110000011011000111110000011001100111101111110100101000101101011000000011100011000111110000101010101010000001000000111010001011011100010110011011111011010000100000111101011000001101001001000000000111110000000100010110111101111101000110010100100000111110011111000101011010111010011011000000101111010001001001100000000000101001010000100000000010000100000111101010111011111001111110011000001100010011001010000001010111101100101111101010001001101010110010011001010101100100111010101001111001101010001011101110010101111110110100000000000111011001000000111001111010001101000110001111100010010111111010010000111000011001110011100111010000111010100100000101100111000010010110100000111001101100110110010011101111111011111111111011001100110101010110001101010000000110110111110100000001001110000111101001000010000111001100000100001110000111011011011000010001101100100000000111111000011000001101000001010111101110101101010000000000110011010100100100100010101010110000010000011011000011111001101000001000101111111101100000111010011110001111100101010000011011101011100011011100100111011011001010000101100101011001011111100011110011101000001110000000111110011010000100100100000000011000111000100001100001001110101010011111101100111101000011010000010101000000001100111000111111011101110001110010001011001100000010011111101110010000101101010110011000100000010000101110011000100001110010010011010100111111011111000010010010111111001111111111000111101000010001101100111010010100010100100001001101001100011000100010110001100100101110000000001110000011111110111010001111100110001001110111001000011011001001110010111100001010111101101110001100101110100000011100010010101110111100101010110111111110001011010111110101010010110011001111111101001101011100110000010001011100101011111110010000000000000110100100011110011110011111000001011000000000011111111111000000000110110000000111111110101100110001000000111000011110000000001001110010110011111000011000000100100010111000000100001111110000110010011001100010010000100100011000010111111111111011111100010111111111100011010100011001101011111101111101011011001011000001101000111000111011101000010100010011000001000011000111111001001110000110010010100110100110110011010110011001111110100100011001110001111100001000100111111001001100011111101100111000101000001100110110110011111100000101111011010011000000100000110110110011111101110101100101001001011110100000100000100000000111110111011001011110001101100000010011100101100001101111001110000111111000101100000001010001010011011001010011110000001011000000001110001111111000110011000011110101011001110010011011001001011011010011101100010000101011001010100011000100000000101110111000110110111001100001111111001110101110101000110010000011010001101011011111000001110011100111100110010001101001110110010001100011111001001010011111000011111101011001001011100010010000000110011001000000000100111011101100101111001001000110101100011000010110010011101001111101001000010100111000111001001111111000111101111000100100010001111101110000100011000010111111000100101011001111110111000000100010101101011100011111111110011000000101111011100000100001101101011110110100100110101101101001101000011000001000011001101101000111100000001111101100000000111011000101000100100001100001101001101001101110111100100100000000010101100110110111111111000001110111100011001000010101111111001110010010111001101101110111001000101100001000110010111001000010100001011100101110110100001011100001110000111001110000000101000000101110011101101111100000110101010001000011010000110001010101001010011100001101101010001111101101000001001101111010000101101101111000011111001110111111001110000100100010110011111011101111000111110110011011101010111000000011100111000000110000011000111010011001101000011101001011010110101110111101101110110010111110111101110111101100001100001000011111111100000010101100111100000011000101001100110110110100110010001010110000100011100011101100000001011010111111110111010010000110000100111110010010111000111011110000110100110000111000010110110000101111110011010111000110111011101000010001010001111111001011011110000011101101110000110011101000101011011010001001000111110111000010000100010111001000001001111101100001111000111001111100001000101100000111011110100111100101111111010101111111011000000001110110001000010001110000101100101111101010000011001100000111001010110000111011010110100101110110111011001100001100100000000010010010101001000111011000000100010011000000100110111111100001011110000001101001100001011001100100010100000001110100110110110011001000111110111111010111100000001111111111101110010001100000110110011100001100101001001111100100111100101101001001110111110101111111100111111101010111000011010100110111001011001111101111000010011100011100010101111000110101110001101000011001001110001001110011010000010010111011100101111001110001001110111110100000111011110000111011000000000010000110101101000111100110000111111110000000011111011000111001000000000101010110001110000001110111111101011010000010111111011100100111011101110001101001001111000100010010010011001110001001101100111010000010001100010100111100011001001110001110011011111111100100110111010100011001111011101111010000110100100110110101010001000010110100000011000100111100100000001011101011110010101100101110110001111010000000110001111111110001000111111011001101100010001001001000001011011000010000100110111001000001101100011000100011000001110111100010111100100001010111010000011001111100111111101100001000110000001000110111111100111000010011110100111100001000111110101000001000000010111110011001111100010111111001000010000011111110111100100101111111011011101100010000110101011011001111000000100110101101111101110110111001011100100111011010001000011111000001101111101010001110001101100000101011000100010111011100001100110010000011110011101110000000100101000111101000111010000011111001000111110000100010001001000001000010011100000111001110001100001011100100000001001001010011001110100000101011100111111011011000000000000001000001101110011110011100001100011101100110111101000101011110111110101100100011110111010000010011111000111000001111000001110001111010001001011101000000101011000001110000001101000001001001100101110101010100000011001011111110010010110000110001010001111001101001100011111001110011010011000001110111000010000011110100110101100001010000001100001110000001111101001111001101011110011000001000100000100001000000001111100111011111010101100111000101110;
localparam PROTOTYPE_DOWN = 10000'b0111000110111000010001010011101111100111000001111111100100110100101111010100000011101010100010111000110001111010111000110101110011011110000001011100000110001111000111100010100010110110000110010111110001111101101111101100010000101011010001111110001110010001110011110000111100001010011100001000100000000001101100001100111101000011100000110110011100101111101010000010000001001110011011100000100100110110011100111001001101000000100000011000000010011010100000011101011100101000110101011011100010000010110010111111001000100000100111110110011011001110100010111110001101110010101000001101110011000111100011011000101101000101101010011111100010100101111010001111011110010111100010100011010101111101100000001001000100111101011011110000111101100110011100000001011100101111110011111110000000011111011101110110000110000111100010100010111101110101111110111111010111100100110011001110000001100011001111100111001110011100000111001001100111001100010111010011000011000111000111101111110110001100001011010100101100100000101001000001110011111001110011100001101111111011000000100000110010110000111101110011000011110111111000011111110101100100011000011101000110111001101010001100010000101111101110111011110001010000110111100000011010100110001110111111010101000111110010111100001111000001100000000010010001000001001111111110010101100100000111011010000000010111110001011000001011111111101100101010111010100101110010010000010101111100101010010010101111000111110011000111111001100100111101001000100001101100010101100110000010100010111110011100001000110001000001100010010010111000111000101001111101100001011101101011100100000100000011010110000111001100011000011110011101000100100101000111011000100110111111111110111111110111011110000110000111010100110110000100011111001100111000011111110100001111101000111110100101110001010011010110011100000110000011110011111110101111110100110100100001000100011100001101001111100111111001100011101111111110010100110111111111000110010000001100111111011110110000000110101101011100010001100000110010000001111100110111101010100111000100110010001101011010101101011110110101010001010110101101000101001010000111000000010011111001111011011001100010100000101110000000011111110001100001000101011000000100110000000110110000001001111011100110001100011111011010111010010111011101110110110110110100010011110001010011101000101010110000010110110010001010000101111001100000001101101000011110000000100100000011110011110000111110101001110011100001011111011010011010000100100001000000101000100110010000001111100100001110110000000011000111011110010010100100000011111001000100011001011101100011110000101100111000011011100010001000000001100001001111101111100110010001011111101000010010010010111011111100000111100101111111101110111001010111010001111100011110110011100000001001111100000111010000100111111110010111000000011111000101001011000111011111000111111000101010000001101111100010011000000001010001010100011011101000001110100111100101101101101100100111111000110001001010011110110101001100010111101110001101000011001111000000100111101111111111011001100001010010101000000001101100101010010101000010011100111111011100110111101100110011010001101000111111110100000001100011110100001001011000001001111011010110001001111110000101001100110111101111000001101010010011101111000000110100001000010101001101111011110001000101010110011011100010011001000111111001001000000001110000111001000101100011011111110010100011001110011000110011110101010100111111101100100100010010001001111110010101100001001111111000001101011100000000000001010010100001011011000010100010101100000010101100001001111011110000001111011100111001010100001011001000001100000011111010011111001011111000110001111101001100111101011001100001000101101011100000000000011000111111100101011110010000101010100100011001111010000001000011111111011000000110000111110001100000011010011000001100111110001100100000110111101111111000110010100100000111110011111011011010001111011011011011000100000110001000001100111111001011000010000100000000010110101001001011010110011100111101110001010001100010011001010000000011011101111010111100110010000100011110011010110100000011101000100111100011000001010000001111110010101000010110111100011010111010001000000111101010111100001000110000111100010010110101110000000100111011001010011100100111000111010100100000001101111000010010110100000111000001101010110010001101111001010010000111011010110111101010100001011000000000111111000010110000011101110100111101110111101111000011100011010001110000111011011011000010000000100110000000000111000000110001101000101010111101110111011010000000000101100000100100100110010010000011100011001101010110011100001101110000111011111111101100101111001000011111000000010010110011101101111000100111100000111011010010000000110111010011111011110100011110000001000001110000100011111001010000100101001101001011000111000000010010001001110101010011101011100110011000001010001110011000001000010011000111111111110000001111001111011111100000010101100010010001100111100000110011001100000010000101110101010111001110010010011010100111111011111000110010110111111001111100111000011101000010001101101111010010100010100010001001101000011101000100010101100000000101110000000011110000010110110111000011111100100001110010110000111101001010000010010111100001010111011101111110000000111000000011101101000100110110100110010110100111111001011010111110101010001001010001111111110001111101100001100010001001100001011111110010000010000000111100100011110011110011111000110011000000000011001110010000000000110110000001011111110101101001101000001111000101110111110011001110011011011111010100000100100000011111001001100101011110000000010000110100010010001000110111000000111111111011011111100010000111111111001010100111001101111111000001101011011100000100000011111111000001011101011110111100000000101000011000101111001110111000101001001010011101001000011010110011011111100001000100001110000111100010101100010011001001000001000101100011100101011111100110110110011111100011010110111101101100101100010110110110011110001110101100100111010011110110000100000000000000011100111101011011110000100111000011011011110100001101010000001100110111100111100011101001111010110111111110111110110001100001110000010001111111000110011000011110100011001110010011011100001011000010001101100011110111011001000100111000001111101001111000000110111000101111011111111001001101111111100101010000111010111100011101111111101110011010111100100011001100111110110110001100011100001111010011010000011111111011001011011100010000001000110101011000000101000111011100100010000101101000110100100011000101000001010101010001101101000100010111000110001001111111000100001111000100101100110011101001111101011000010111111110000101010101111110011000000100011101101011100011111111110010000000100000111100011100001110001011110110110100110100111100111101010011000001001111001111101000111100000000111001101000011010101100100100110100001100001101001101001111111000100111111000000010110000111011000000101111111001001100011001000111010000111111111110100001001101101110101110010001001101000110010111001000110000011011100101000000100111000100011100000111001110100000101000011110110000100001100100110010101110001000011010000110001010101001010011100001101101010001001101101000000111110011010111001101001111000011111001110111111010010100100100100110101011111101111000100011110100111011101110000000011100111000000110000000000000010011001101101110110101110000101001111111011110110110100111110111101110100001100101100110000011111101101000010111011011100000011000100001100110110110100110010011010010000100010100011101100000001010110111100000011000010011101000000111111010010111111111011110000110100101110111000010010100000001001010011010111100010011011101011010111110001111110110011000110000011111011110000000011101000101011001011101000011111001111011010000100010111001001001001011101110100011100111001111100100011101100000111011110100111100011110000101001001110101101110001111010001100010001110100101100101101101100000011001100000110101100111111011011101001100001110110110011001101101100100000010011110010101001000010100110100110001111011100100110100011100111101110011101101001101110011101100011110100000001110100011000110011000000011010010011010110000001100001111011011110010001110000110001011100001100100001101111010110001100110011001001010111111001111100101111111101010111000011010000010000001000101111101111000010000010000010010001011111110000010110001000011010110001000111100011011111110000111011110001100101110001001110011110100000111011001111010011000000000010000110101101000111100110000111111110000000011111000100100010110000001101010111011101101001110011100111001000000010111111011101100011011110110001100001001110100110010010011011100000001011111100110010001010001100010101101000011001000110110110011011011110101100111110010011011001111011101011100001010000100110110101010001010010110100001100100000111110000000001011110110011010111100101001001111110010000000110001111100100001010011111010001101100010001011001000001011000000110000100110100111000001100100111110100000111011110100101101000100000001010111011110011101111100111000101111100111110000001000000011110100111000010011111100100000110110111100001111110000000001000011110000011100010011111001000010110011111000000100111001111111011011101101110000110111000000100111000010000110101101111101010001111000000100111111011010001000010110000101101111100000001011101101100000111011001010010000111011001110111100000010110000101110000001000101000111101010101001000000001001100111111000000000001001000001110010001000010001111110001010001011001111000101001101010101010010100001101101100111111011100110001000000001000110000001100000011001110011111001100110111110100111101110111110101101100011110111010000010011111000111000000110100000100111110010101101011101000000110011000111100110001101000000111011100011000101010100010100110010001110010010110000010001000110011001110001101111111011111100010011000001110111000010000001110111111101001001010000001100000010000001111101001111001101011110011000011011111100110001000000001111100010001111010000110100000101110;

    hv_binary_adder #(
        .AM_NUM_FOLDS       (AM_FOLD_WIDTH),
        .AM_NUM_FOLDS_WIDTH (AM_NUM_FOLDS_WIDTH),
        .AM_FOLD_WIDTH      (AM_FOLD_WIDTH)
    ) BIN_ADDER (
        .hv         (similarity_hv),
        .distance   (distance)
    );

    assign hvin_fire    = hvin_valid && hvin_ready;
    assign hvin_ready   = prototype_counter == 0 && fold_counter == 0;

    assign dout_fire    = dout_valid && dout_ready;
    assign dout_valid   = prototype_counter == 10;

    always @(posedge clk) begin
        if (rst || dout_fire)
            prototype_counter   <= 0;
        else if (fold_counter == AM_NUM_FOLDS-1)
            prototype_counter   <= prototype_counter + 1;
    end

    always @(posedge clk) begin
        if (rst || fold_counter == AM_NUM_FOLDS-1 || dout_fire)
            fold_counter    <= 0;
        else if (hvin_fire || (fold_counter > 0 && fold_counter < AM_NUM_FOLDS-1) ||
                        (fold_counter == 0 && prototype_counter > 0 && prototype_counter < 10))
            fold_counter    <= fold_counter + 1;
    end

    always @(*) begin
        case (prototype_counter)
            0: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_ON[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            1: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_OFF[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            2: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_GO[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            3: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_STOP[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            4: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_LEFT[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            5: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_RIGHT[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            6: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_YES[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            7: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_NO[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            8: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_UP[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            9: similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_DOWN[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
            default: similarity_hv = {AM_FOLD_WIDTH{1'b0}};
        endcase
    end

    always @(posedge clk) begin
        if (prototype_counter == 0)
            distance_ON <= (fold_counter == 0) ? distance : distance_ON + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 1)
            distance_OFF <= (fold_counter == 0) ? distance : distance_OFF + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 2)
            distance_GO <= (fold_counter == 0) ? distance : distance_GO + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 3)
            distance_STOP <= (fold_counter == 0) ? distance : distance_STOP + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 4)
            distance_LEFT <= (fold_counter == 0) ? distance : distance_LEFT + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 5)
            distance_RIGHT <= (fold_counter == 0) ? distance : distance_RIGHT + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 6)
            distance_YES <= (fold_counter == 0) ? distance : distance_YES + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 7)
            distance_NO <= (fold_counter == 0) ? distance : distance_NO + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 8)
            distance_UP <= (fold_counter == 0) ? distance : distance_UP + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 9)
            distance_DOWN <= (fold_counter == 0) ? distance : distance_DOWN + distance;
    end

    always @(posedge clk) begin
        if (prototype_counter == 1 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_OFF + distance < distance_ON) ? 1 : 0;
            curr_min    <= (distance_OFF + distance < distance_ON) ? distance_OFF + distance : distance_ON;
        end else if (prototype_counter == 2 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_GO + distance < curr_min) ? 2 : keyword;
            curr_min    <= (distance_GO + distance < curr_min) ? distance_GO + distance : curr_min;
        end else if (prototype_counter == 3 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_STOP + distance < curr_min) ? 3 : keyword;
            curr_min    <= (distance_STOP + distance < curr_min) ? distance_STOP + distance : curr_min;
        end else if (prototype_counter == 4 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_LEFT + distance < curr_min) ? 4 : keyword;
            curr_min    <= (distance_LEFT + distance < curr_min) ? distance_LEFT + distance : curr_min;
        end else if (prototype_counter == 5 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_RIGHT + distance < curr_min) ? 5 : keyword;
            curr_min    <= (distance_RIGHT + distance < curr_min) ? distance_RIGHT + distance : curr_min;
        end else if (prototype_counter == 6 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_YES + distance < curr_min) ? 6 : keyword;
            curr_min    <= (distance_YES + distance < curr_min) ? distance_YES + distance : curr_min;
        end else if (prototype_counter == 7 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_NO + distance < curr_min) ? 7 : keyword;
            curr_min    <= (distance_NO + distance < curr_min) ? distance_NO + distance : curr_min;
        end else if (prototype_counter == 8 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_UP + distance < curr_min) ? 8 : keyword;
            curr_min    <= (distance_UP + distance < curr_min) ? distance_UP + distance : curr_min;
        end else if (prototype_counter == 9 && fold_counter == AM_NUM_FOLDS-1) begin
            keyword     <= (distance_DOWN + distance < curr_min) ? 9 : keyword;
            curr_min    <= (distance_DOWN + distance < curr_min) ? distance_DOWN + distance : curr_min;
        end
    end

endmodule : associative_memory
